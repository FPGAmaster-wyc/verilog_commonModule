library verilog;
use verilog.vl_types.all;
entity key_filter_tb is
end key_filter_tb;
