library verilog;
use verilog.vl_types.all;
entity page_rd_tb is
end page_rd_tb;
