library verilog;
use verilog.vl_types.all;
entity edge_detection_tb is
end edge_detection_tb;
