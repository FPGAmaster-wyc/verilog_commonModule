library verilog;
use verilog.vl_types.all;
entity freq_ji_tb is
end freq_ji_tb;
