begin
	$[![]!]
end



case ($[![]!])

endcase



always @ (posedge clk)
begin
	if(!rst_n)
		begin
			$[![]!]
		end	
	else
		begin
		
		end 
end 

else if ($[![]!])
	begin
	
	end 

/*    */