library verilog;
use verilog.vl_types.all;
entity page_wr_tb is
end page_wr_tb;
