library verilog;
use verilog.vl_types.all;
entity key_scan_tb is
end key_scan_tb;
